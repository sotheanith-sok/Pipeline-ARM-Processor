`timescale 1ns / 1ps
module IM(in, out);
	input 	[63:0] in;
	output	[31:0] out;



endmodule
