`timescale 1ns / 1ps
module InstructionMemory(Address, out);
	input		[63:0] Address;
	output [31:0] out;
	
	reg	[7:0] IM	[0:225];
	
	assign out={IM[Address+0], IM[Address+1], IM[Address+2], IM[Address+3]};
	
	initial 
		begin
			//LDUR X1, [X31, # 8]	
			{IM[0],IM[1],IM[2],IM[3]}=	32'b11111000010_000001000_00_11111_00001;
			//LDUR X2, [X31, # 16]	
			{IM[4],IM[5],IM[6],IM[7]}=	32'b11111000010_000010000_00_11111_00010;
			//LDUR X3, [X31, # 24]	
			{IM[8],IM[9],IM[10],IM[11]}=	32'b11111000010_000011000_00_11111_00011;
			//LDUR X4, [X31, # 32]	
			{IM[12],IM[13],IM[14],IM[15]}=32'b11111000010_000100000_00_11111_00100;
			//LDUR X5, [X31, # 40]	
			{IM[16],IM[17],IM[18],IM[19]}=32'b11111000010_000101000_00_11111_00101;
			//LDUR X6, [X31, # 48]	
			{IM[20],IM[21],IM[22],IM[23]}=32'b11111000010_000110000_00_11111_00110;
			//LDUR X7, [X31, # 56]	
			{IM[24],IM[25],IM[26],IM[27]}=32'b11111000010_000111000_00_11111_00111;
			//LDUR X8, [X31, # 64]	
			{IM[28],IM[29],IM[30],IM[31]}=32'b11111000010_001000000_00_11111_01000;
			//LDUR X9, [X31, # 72]	
			{IM[32],IM[33],IM[34],IM[35]}=32'b11111000010_001001000_00_11111_01001;
			//LDUR X10, [X31, # 80]	
			{IM[36],IM[37],IM[38],IM[39]}=32'b11111000010_001010000_00_11111_01010;
			//LDUR X11, [X31, # 88]	
			{IM[40],IM[41],IM[42],IM[43]}=32'b11111000010_001011000_00_11111_01011;
			//LDUR X12, [X31, # 96]	
			{IM[44],IM[45],IM[46],IM[47]}=32'b11111000010_001100000_00_11111_01100;
			//ADD X2, X1, X3
			{IM[48],IM[49],IM[50],IM[51]}=32'b10001011000_00011_000000_00001_00010;
			//SUB X6, X5, X4
			{IM[52],IM[53],IM[54],IM[55]}=32'b11001011000_00100_000000_00101_00110;
			//OR X9, X7, X8
			{IM[56],IM[57],IM[58],IM[59]}=32'b10101010000_01000_000000_00111_01001;
			//AND X12, X10, X11
			{IM[60],IM[61],IM[62],IM[63]}=32'b10001010000_01011_000000_01010_01100;
			
			
		end
endmodule
